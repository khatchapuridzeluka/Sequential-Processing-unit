module au (
	input [31:0] a,
	input [31:0] b,
	input u,
	input sub,
	output [31:0] s,
	output neg,
	output ovf
);

 

endmodule 