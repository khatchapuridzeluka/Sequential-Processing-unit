module instruction_decod_helper (
	input [31:0] instruction;
);


endmodule 