module instruction_exe (
	input clk,
	input [31:0] instruction,
	output t
);

endmodule 