module alu(
	input [2:0] optype;
	input [4:0] rs;
	input [4:0] rt;
	input [4:0] rd;
	
);

endmodule 